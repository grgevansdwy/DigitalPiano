module encoder(in, out);
	input logic [4:0] in;
	output logic [31:0] out;
	
endmodule	